PK   0g}T]D�@  a�     cirkitFile.json�]Yo�8�+ͫe��a�mg�f��^�>$�@[TGXG��r��Rr�K�J܃M#I۬���X,�h�W�/�L7�J�_t�/v�w�Åw���z�.[xwE�ֻ�s��n����_�����*[�O�ĉZ%���(�~�$�����_+�9�D�K�?�������ە��SF	c��D�~���Q�ϕ��阇z�Jo1�1h��&�(?���:1$�&�!_�u�b�7�y�!�C���`�jN��,�Hh&� 1�׋�'͛�� G����n�㾠��~��~H�F`F�XXf$��E`i��E`i��E`i��E`�
������`0����!6�q<��K4���K4��L4���L4�����L�?�&�����<�.;�ۜ�q�'���3�9��un�{����_]��+Z�j�x�W��9$F���9�)[l��H����Q�#U/���X-�іczO�3���H���R�)|�>�V��9)|��D
_b��t%R��-]�໻X�z���M�N��5�������T�CsԡݳX~��V�nsEI`)=M��'lv�]������X���y�zV���/PS��~��D�ǈS14@�
�)��0"j
�4����r9#"��xNÈ�)��0"j
�4����2;#"���NC�
�-�q"�ۜ,pS!��y"Nd���o*��tOĉ,~s� �B�^�'@q̷�E~9��N/�pq�fz	� ű�N/��8ֱ�}
��������a��4��S��Q0Q��4捈��1�004*4*D1X�_;Ϩ�S��Q��Q��Q��Q�X�#�C��X	.�S��4*�4*�D���%���IC��(�����˹�|��D�V�_^�E�{Z�~�_�E�3	h��q��
��Z՚�p\�C]�-�pL ��I��cFD@mᘄP[8&aD��I��cFD@mᘄP[8&aD��I�4!�.jӅm����7ұpLÉ,vs��M�t,�p"�ߜ,���f��(��6�p�GqhzF����͌�1ű��(�Q�؜�1�z]~N� �F���7�pL C�aN#bN�bA�bA�iT,hT,hT,hT,hT,hT,hT,hT,iT,iT,�R	K˓*��('�	\8ƣ�%p��r�_��c<
M�<�����[��7N��w�Zx_�J�ӻ���,-�tWe��..���1�p�8���9.��<P�{�G��L�q����0��g�u��ó�]Љ}�'f�#4�R�1π?��ϝ���l��>���a�����Y�T���{���9�k{�sr?y�pV���r�?�ġ��7�NH4�MR^�7�U�+vZo�6����юx���z��'tx���5#4���6�;{�n�=�����q����]�{���EF������{�R�.�'T�m��!I	,�C���,��9$4D�I��n�C�@C���,��8$4D���q�膤��8nn�� ��� ��1��ذ<b('�x��f5,�8�	�cƦ4��`��؈��'ҹ{�0t�����?X�f�9����9��P XA#�]e=E�?��"�%:�p�,�md�>E��:X�
t�'��l#C��T`u*�:X����?j�Z�:�X�J�
���
S� L�>0����Ќ�`��	�'�y��0X��s�=x����`�x��@��	��l����m��w��L{����@Z�Y�����wl��m1�Ak�ZKnM���֘[kn͹��ց[a=D�m=���CXa=��h�	�!�����c=���v����#�����>��vl�kۯi�d��4�=��Mj([��_1�i�p�۷4�&���#�2�+�ᴘ�Y�p�|`�{�iB�v��V����������_�$���ib�&~l��&yl�æ���x�����6�2ߥ�b_�>ˢ<
E���Y����O2��<_m�z���H�"�Wu��L�:�m�b�������I���Xz����Gz�ǡ��M����h��P��tU�Y�n�J��j��ᾮ��9�R��׶u�}Qۃ}������s(��3���쾾/�jp���r2�{]}*��z�߫�E�3�6�j�V��\m�C���<7{Ƥ��I��>sd�/��/a^�<��aGt���e�\��k-�w��'�2�b��zf���X�a�1��U$vi2E��M��+ޮ*�ة��g�ԌhQm��8��l"�d����x��{�v��� ^ċCWK�:���|";j$����g�=�p�%!�.�-�瑖�q����q����8��$�sz瑖�q��N��y���3:�#v��<�{g9h	V�2���μ����0�������n�h�)��!+v�� �Ǘ|��R�]�V���L�ա�yWf�cN�z��<Z���L����J�*Ʉ`fx֙YnV�߬��gIq�%׬�X����Fb6�yp!�d��7$=��y���cr)�" _D�-d-����p���r_�̏$0rHb&�Wb�Z�,ֲ/!P� ��dH1ib�X	W��i[B���9%7���e�Ȭ��5
[$s2�uą�ˇ�׳����fh��ݍ.>�X�p/W�7��=�w�mKmnt���ŇJ���O���o��{u���k>!y�]\=<���[\���P�ﲦi~�A�e�"�(�@U��GRn��t��vEYP�M�����ʳWr����c3���݋K��������Z,�ޑ9�*�٘U'��uC�~}���u��>@�E�̨��+��R�;X�v�,��'@M�NUS�6>>�&Y�L0�,�d�Of�#�Y���A{���tʃa_Sy�4��yq������1�����b3���V�M�q��&P�*:CD' r�e�P39X�ǥ�>�2���
vW�8����j=df�Zp�Vq�PZ7&͠j�Mn8����7�]M��̮�גޥ"��O �}��x͙@��F��v��i�ӭ��������J��S�"sb�T8�z�!��=��9�ث9�\����9��[}��C\��83�C	�:ԫ[B�\K�-Z����wU�P۽wa��o^����<��o��w���[�����PK
   0g}T]D�@  a�                   cirkitFile.jsonPK      =   m    